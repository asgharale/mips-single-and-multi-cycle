module InstrMemory (
    input [31:0] PC, 
    output [31:0] Instr
);
    reg [31:0] mem [0:255];

    initial begin
        mem[0] = 32'b00000000000000010000000000100000;
        mem[1] = 32'b10001100000000010000000000000100;
        mem[2] = 32'b10101100001000100000000000000000;
        mem[3] = 32'b00010000001000100000000000000100;
        mem[4] = 32'b00001000000000000000000000000000;
    end

    assign Instr = mem[PC >> 2];
endmodule